// ADCinterface_qsys.v

// Generated using ACDS version 14.1 186 at 2015.05.23.22:54:30

`timescale 1 ps / 1 ps
module ADCinterface_qsys (
		input  wire [7:0] adc_dataandclock_adc_data, //   adc_dataandclock.adc_data
		input  wire       adc_dataandclock_adc_clk,  //                   .adc_clk
		output wire       adc_interface_adc_csbn,    //      adc_interface.adc_csbn
		output wire       adc_interface_adc_sdio,    //                   .adc_sdio
		output wire       adc_interface_adc_sclk,    //                   .adc_sclk
		output wire       adc_interface_adc_oen,     //                   .adc_oen
		output wire       adc_interface_adc_sdon,    //                   .adc_sdon
		output wire       adc_interface_cha_3p5,     //                   .cha_3p5
		output wire       adc_interface_cha_2x,      //                   .cha_2x
		output wire       adc_interface_cha_8p5x,    //                   .cha_8p5x
		output wire       adc_interface_cha_in1,     //                   .cha_in1
		output wire       adc_interface_cha_in3,     //                   .cha_in3
		output wire       adc_interface_cha_en,      //                   .cha_en
		output wire       adc_interface_cha_in4,     //                   .cha_in4
		output wire       adc_interface_mon_fs,      //                   .mon_fs
		output wire       adc_interface_mon_en,      //                   .mon_en
		output wire       adc_interface_chb_en,      //                   .chb_en
		output wire       adc_interface_chb_in2,     //                   .chb_in2
		output wire       adc_interface_chb_in1,     //                   .chb_in1
		output wire       adc_interface_chb_in4,     //                   .chb_in4
		output wire       adc_interface_chb_3p5x,    //                   .chb_3p5x
		output wire       adc_interface_chb_2x,      //                   .chb_2x
		output wire       adc_interface_chb_8p5x,    //                   .chb_8p5x
		input  wire       buttonsandswitches_b1,     // buttonsandswitches.b1
		input  wire       buttonsandswitches_b2,     //                   .b2
		input  wire       buttonsandswitches_sw1,    //                   .sw1
		input  wire       buttonsandswitches_sw2,    //                   .sw2
		input  wire       buttonsandswitches_sw3,    //                   .sw3
		input  wire       clk_clk,                   //                clk.clk
		output wire [7:0] leds_led                   //               leds.led
	);

	wire         master_0_master_reset_reset;                               // master_0:master_reset_reset -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_001:reset_in1]
	wire  [31:0] master_0_master_readdata;                                  // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                               // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                   // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                      // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                             // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                     // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                 // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire   [7:0] mm_interconnect_0_adcinterface_0_avalon_slave_0_readdata;  // ADCinterface_0:readdata -> mm_interconnect_0:ADCinterface_0_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_0_adcinterface_0_avalon_slave_0_address;   // mm_interconnect_0:ADCinterface_0_avalon_slave_0_address -> ADCinterface_0:address
	wire         mm_interconnect_0_adcinterface_0_avalon_slave_0_read;      // mm_interconnect_0:ADCinterface_0_avalon_slave_0_read -> ADCinterface_0:read
	wire         mm_interconnect_0_adcinterface_0_avalon_slave_0_write;     // mm_interconnect_0:ADCinterface_0_avalon_slave_0_write -> ADCinterface_0:write
	wire   [7:0] mm_interconnect_0_adcinterface_0_avalon_slave_0_writedata; // mm_interconnect_0:ADCinterface_0_avalon_slave_0_writedata -> ADCinterface_0:writedata
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [ADCinterface_0:rst, mm_interconnect_0:ADCinterface_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> master_0:clk_reset_reset

	ADCinterface adcinterface_0 (
		.read         (mm_interconnect_0_adcinterface_0_avalon_slave_0_read),      //     avalon_slave_0.read
		.write        (mm_interconnect_0_adcinterface_0_avalon_slave_0_write),     //                   .write
		.readdata     (mm_interconnect_0_adcinterface_0_avalon_slave_0_readdata),  //                   .readdata
		.address      (mm_interconnect_0_adcinterface_0_avalon_slave_0_address),   //                   .address
		.writedata    (mm_interconnect_0_adcinterface_0_avalon_slave_0_writedata), //                   .writedata
		.main_clk     (clk_clk),                                                   //         clock_sink.clk
		.rst          (rst_controller_reset_out_reset),                            //         reset_sink.reset
		.ADC_CSBn     (adc_interface_adc_csbn),                                    //      ADC_Interface.adc_csbn
		.ADC_SDIO     (adc_interface_adc_sdio),                                    //                   .adc_sdio
		.ADC_SCLK     (adc_interface_adc_sclk),                                    //                   .adc_sclk
		.ADC_OEn      (adc_interface_adc_oen),                                     //                   .adc_oen
		.ADC_SDOn     (adc_interface_adc_sdon),                                    //                   .adc_sdon
		.CHA_3P5X_PDn (adc_interface_cha_3p5),                                     //                   .cha_3p5
		.CHA_2X_PDn   (adc_interface_cha_2x),                                      //                   .cha_2x
		.CHA_8P5X_PDn (adc_interface_cha_8p5x),                                    //                   .cha_8p5x
		.CHA_IN1      (adc_interface_cha_in1),                                     //                   .cha_in1
		.CHA_IN3      (adc_interface_cha_in3),                                     //                   .cha_in3
		.CHA_EN       (adc_interface_cha_en),                                      //                   .cha_en
		.CHA_IN4      (adc_interface_cha_in4),                                     //                   .cha_in4
		.MON_FS       (adc_interface_mon_fs),                                      //                   .mon_fs
		.MON_EN       (adc_interface_mon_en),                                      //                   .mon_en
		.CHB_EN       (adc_interface_chb_en),                                      //                   .chb_en
		.CHB_IN2      (adc_interface_chb_in2),                                     //                   .chb_in2
		.CHB_IN1      (adc_interface_chb_in1),                                     //                   .chb_in1
		.CHB_IN4      (adc_interface_chb_in4),                                     //                   .chb_in4
		.CHB_3P5X_PDn (adc_interface_chb_3p5x),                                    //                   .chb_3p5x
		.CHB_2X_PDn   (adc_interface_chb_2x),                                      //                   .chb_2x
		.CHB_8P5X_PDn (adc_interface_chb_8p5x),                                    //                   .chb_8p5x
		.D            (adc_dataandclock_adc_data),                                 //   ADC_DataAndClock.adc_data
		.DCO          (adc_dataandclock_adc_clk),                                  //                   .adc_clk
		.button1      (buttonsandswitches_b1),                                     // ButtonsAndSwitches.b1
		.button2      (buttonsandswitches_b2),                                     //                   .b2
		.switch1      (buttonsandswitches_sw1),                                    //                   .sw1
		.switch2      (buttonsandswitches_sw2),                                    //                   .sw2
		.switch3      (buttonsandswitches_sw3),                                    //                   .sw3
		.led          (leds_led)                                                   //               LEDs.led
	);

	ADCinterface_qsys_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                            //          clk.clk
		.clk_reset_reset      (rst_controller_001_reset_out_reset), //    clk_reset.reset
		.master_address       (master_0_master_address),            //       master.address
		.master_readdata      (master_0_master_readdata),           //             .readdata
		.master_read          (master_0_master_read),               //             .read
		.master_write         (master_0_master_write),              //             .write
		.master_writedata     (master_0_master_writedata),          //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),        //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid),      //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),         //             .byteenable
		.master_reset_reset   (master_0_master_reset_reset)         // master_reset.reset
	);

	ADCinterface_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                         (clk_clk),                                                   //                                       clk_0_clk.clk
		.ADCinterface_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // ADCinterface_0_reset_sink_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                            //        master_0_clk_reset_reset_bridge_in_reset.reset
		.master_0_master_address                               (master_0_master_address),                                   //                                 master_0_master.address
		.master_0_master_waitrequest                           (master_0_master_waitrequest),                               //                                                .waitrequest
		.master_0_master_byteenable                            (master_0_master_byteenable),                                //                                                .byteenable
		.master_0_master_read                                  (master_0_master_read),                                      //                                                .read
		.master_0_master_readdata                              (master_0_master_readdata),                                  //                                                .readdata
		.master_0_master_readdatavalid                         (master_0_master_readdatavalid),                             //                                                .readdatavalid
		.master_0_master_write                                 (master_0_master_write),                                     //                                                .write
		.master_0_master_writedata                             (master_0_master_writedata),                                 //                                                .writedata
		.ADCinterface_0_avalon_slave_0_address                 (mm_interconnect_0_adcinterface_0_avalon_slave_0_address),   //                   ADCinterface_0_avalon_slave_0.address
		.ADCinterface_0_avalon_slave_0_write                   (mm_interconnect_0_adcinterface_0_avalon_slave_0_write),     //                                                .write
		.ADCinterface_0_avalon_slave_0_read                    (mm_interconnect_0_adcinterface_0_avalon_slave_0_read),      //                                                .read
		.ADCinterface_0_avalon_slave_0_readdata                (mm_interconnect_0_adcinterface_0_avalon_slave_0_readdata),  //                                                .readdata
		.ADCinterface_0_avalon_slave_0_writedata               (mm_interconnect_0_adcinterface_0_avalon_slave_0_writedata)  //                                                .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (master_0_master_reset_reset),    // reset_in0.reset
		.reset_in1      (master_0_master_reset_reset),    // reset_in1.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (master_0_master_reset_reset),        // reset_in0.reset
		.reset_in1      (master_0_master_reset_reset),        // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
